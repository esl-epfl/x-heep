// Copyright EPFL contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

module ams_adc_1b (
    input logic [1:0] sel,
    output logic out
);

endmodule : ams_adc_1b

