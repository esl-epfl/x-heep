/*
 * Copyright 2024 EPFL
 * Solderpad Hardware License, Version 2.1, see LICENSE.md for details.
 * SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 *
 * Author: Tommaso Terzano <tommaso.terzano@epfl.ch>
 *                         <tommaso.terzano@gmail.com>
 *  
 * Info: This module defines parameters for the Smart Peripheral Controller extension.
 */

package ao_spc_pkg;

  localparam int AO_SPC_NUM = 1;

endpackage
