/* verilator lint_off DECLFILENAME */

interface if_bundle__pad_ring__root ();
  logic rst_n;
  logic clk;
  logic muxer_pad_connector_pdm2pcm0_pdm_0_i;
  logic muxer_pad_connector_pdm2pcm0_pdm_0_o;
  logic muxer_pad_connector_pdm2pcm0_pdm_0_oe;
  logic muxer_pad_connector_pdm2pcm0_pdm_clk_0_i;
  logic muxer_pad_connector_pdm2pcm0_pdm_clk_0_o;
  logic muxer_pad_connector_pdm2pcm0_pdm_clk_0_oe;
  logic muxer_pad_connector_i2s0_sck_0_i;
  logic muxer_pad_connector_i2s0_sck_0_o;
  logic muxer_pad_connector_i2s0_sck_0_oe;
  logic muxer_pad_connector_i2s0_ws_0_i;
  logic muxer_pad_connector_i2s0_ws_0_o;
  logic muxer_pad_connector_i2s0_ws_0_oe;
  logic muxer_pad_connector_i2s0_sd_0_i;
  logic muxer_pad_connector_i2s0_sd_0_o;
  logic muxer_pad_connector_i2s0_sd_0_oe;
  logic muxer_pad_connector_spi_host1_csb_0_i;
  logic muxer_pad_connector_spi_host1_csb_0_o;
  logic muxer_pad_connector_spi_host1_csb_0_oe;
  logic muxer_pad_connector_spi_host1_csb_1_i;
  logic muxer_pad_connector_spi_host1_csb_1_o;
  logic muxer_pad_connector_spi_host1_csb_1_oe;
  logic muxer_pad_connector_spi_host1_sck_0_i;
  logic muxer_pad_connector_spi_host1_sck_0_o;
  logic muxer_pad_connector_spi_host1_sck_0_oe;
  logic muxer_pad_connector_spi_host1_sd_0_i;
  logic muxer_pad_connector_spi_host1_sd_0_o;
  logic muxer_pad_connector_spi_host1_sd_0_oe;
  logic muxer_pad_connector_spi_host1_sd_1_i;
  logic muxer_pad_connector_spi_host1_sd_1_o;
  logic muxer_pad_connector_spi_host1_sd_1_oe;
  logic muxer_pad_connector_spi_host1_sd_2_i;
  logic muxer_pad_connector_spi_host1_sd_2_o;
  logic muxer_pad_connector_spi_host1_sd_2_oe;
  logic muxer_pad_connector_spi_host1_sd_3_i;
  logic muxer_pad_connector_spi_host1_sd_3_o;
  logic muxer_pad_connector_spi_host1_sd_3_oe;
  logic muxer_pad_connector_i2c0_scl_0_i;
  logic muxer_pad_connector_i2c0_scl_0_o;
  logic muxer_pad_connector_i2c0_scl_0_oe;
  logic muxer_pad_connector_i2c0_sda_0_i;
  logic muxer_pad_connector_i2c0_sda_0_o;
  logic muxer_pad_connector_i2c0_sda_0_oe;
  modport root(
      input rst_n,
      input clk,
      input muxer_pad_connector_pdm2pcm0_pdm_0_i,
      output muxer_pad_connector_pdm2pcm0_pdm_0_o,
      output muxer_pad_connector_pdm2pcm0_pdm_0_oe,
      input muxer_pad_connector_pdm2pcm0_pdm_clk_0_i,
      output muxer_pad_connector_pdm2pcm0_pdm_clk_0_o,
      output muxer_pad_connector_pdm2pcm0_pdm_clk_0_oe,
      input muxer_pad_connector_i2s0_sck_0_i,
      output muxer_pad_connector_i2s0_sck_0_o,
      output muxer_pad_connector_i2s0_sck_0_oe,
      input muxer_pad_connector_i2s0_ws_0_i,
      output muxer_pad_connector_i2s0_ws_0_o,
      output muxer_pad_connector_i2s0_ws_0_oe,
      input muxer_pad_connector_i2s0_sd_0_i,
      output muxer_pad_connector_i2s0_sd_0_o,
      output muxer_pad_connector_i2s0_sd_0_oe,
      input muxer_pad_connector_spi_host1_csb_0_i,
      output muxer_pad_connector_spi_host1_csb_0_o,
      output muxer_pad_connector_spi_host1_csb_0_oe,
      input muxer_pad_connector_spi_host1_csb_1_i,
      output muxer_pad_connector_spi_host1_csb_1_o,
      output muxer_pad_connector_spi_host1_csb_1_oe,
      input muxer_pad_connector_spi_host1_sck_0_i,
      output muxer_pad_connector_spi_host1_sck_0_o,
      output muxer_pad_connector_spi_host1_sck_0_oe,
      input muxer_pad_connector_spi_host1_sd_0_i,
      output muxer_pad_connector_spi_host1_sd_0_o,
      output muxer_pad_connector_spi_host1_sd_0_oe,
      input muxer_pad_connector_spi_host1_sd_1_i,
      output muxer_pad_connector_spi_host1_sd_1_o,
      output muxer_pad_connector_spi_host1_sd_1_oe,
      input muxer_pad_connector_spi_host1_sd_2_i,
      output muxer_pad_connector_spi_host1_sd_2_o,
      output muxer_pad_connector_spi_host1_sd_2_oe,
      input muxer_pad_connector_spi_host1_sd_3_i,
      output muxer_pad_connector_spi_host1_sd_3_o,
      output muxer_pad_connector_spi_host1_sd_3_oe,
      input muxer_pad_connector_i2c0_scl_0_i,
      output muxer_pad_connector_i2c0_scl_0_o,
      output muxer_pad_connector_i2c0_scl_0_oe,
      input muxer_pad_connector_i2c0_sda_0_i,
      output muxer_pad_connector_i2c0_sda_0_o,
      output muxer_pad_connector_i2c0_sda_0_oe
  );
  modport pad_ring(
      output rst_n,
      output clk,
      output muxer_pad_connector_pdm2pcm0_pdm_0_i,
      input muxer_pad_connector_pdm2pcm0_pdm_0_o,
      input muxer_pad_connector_pdm2pcm0_pdm_0_oe,
      output muxer_pad_connector_pdm2pcm0_pdm_clk_0_i,
      input muxer_pad_connector_pdm2pcm0_pdm_clk_0_o,
      input muxer_pad_connector_pdm2pcm0_pdm_clk_0_oe,
      output muxer_pad_connector_i2s0_sck_0_i,
      input muxer_pad_connector_i2s0_sck_0_o,
      input muxer_pad_connector_i2s0_sck_0_oe,
      output muxer_pad_connector_i2s0_ws_0_i,
      input muxer_pad_connector_i2s0_ws_0_o,
      input muxer_pad_connector_i2s0_ws_0_oe,
      output muxer_pad_connector_i2s0_sd_0_i,
      input muxer_pad_connector_i2s0_sd_0_o,
      input muxer_pad_connector_i2s0_sd_0_oe,
      output muxer_pad_connector_spi_host1_csb_0_i,
      input muxer_pad_connector_spi_host1_csb_0_o,
      input muxer_pad_connector_spi_host1_csb_0_oe,
      output muxer_pad_connector_spi_host1_csb_1_i,
      input muxer_pad_connector_spi_host1_csb_1_o,
      input muxer_pad_connector_spi_host1_csb_1_oe,
      output muxer_pad_connector_spi_host1_sck_0_i,
      input muxer_pad_connector_spi_host1_sck_0_o,
      input muxer_pad_connector_spi_host1_sck_0_oe,
      output muxer_pad_connector_spi_host1_sd_0_i,
      input muxer_pad_connector_spi_host1_sd_0_o,
      input muxer_pad_connector_spi_host1_sd_0_oe,
      output muxer_pad_connector_spi_host1_sd_1_i,
      input muxer_pad_connector_spi_host1_sd_1_o,
      input muxer_pad_connector_spi_host1_sd_1_oe,
      output muxer_pad_connector_spi_host1_sd_2_i,
      input muxer_pad_connector_spi_host1_sd_2_o,
      input muxer_pad_connector_spi_host1_sd_2_oe,
      output muxer_pad_connector_spi_host1_sd_3_i,
      input muxer_pad_connector_spi_host1_sd_3_o,
      input muxer_pad_connector_spi_host1_sd_3_oe,
      output muxer_pad_connector_i2c0_scl_0_i,
      input muxer_pad_connector_i2c0_scl_0_o,
      input muxer_pad_connector_i2c0_scl_0_oe,
      output muxer_pad_connector_i2c0_sda_0_i,
      input muxer_pad_connector_i2c0_sda_0_o,
      input muxer_pad_connector_i2c0_sda_0_oe
  );
endinterface

interface if_bundle__core_v_mini_mcu__pad_ring ();
  logic jtag_tck;
  logic jtag_tms;
  logic jtag_trst_n;
  logic jtag_tdi;
  logic jtag_tdo;
  modport core_v_mini_mcu(
      input jtag_tck,
      input jtag_tms,
      input jtag_trst_n,
      input jtag_tdi,
      output jtag_tdo
  );
  modport pad_ring(
      output jtag_tck,
      output jtag_tms,
      output jtag_trst_n,
      output jtag_tdi,
      input jtag_tdo
  );
endinterface

interface if_bundle__ao_periph__pad_ring ();
  logic boot_select;
  logic execute_from_flash;
  logic exit_valid;
  logic spi_flash_sck_o;
  logic spi_flash_sck_en_o;
  logic spi_flash_csb_0_o;
  logic spi_flash_csb_0_en_o;
  logic spi_flash_csb_1_o;
  logic spi_flash_csb_1_en_o;
  logic spi_flash_sd_0_o;
  logic spi_flash_sd_0_en_o;
  logic spi_flash_sd_0_i;
  logic spi_flash_sd_1_o;
  logic spi_flash_sd_1_en_o;
  logic spi_flash_sd_1_i;
  logic spi_flash_sd_2_o;
  logic spi_flash_sd_2_en_o;
  logic spi_flash_sd_2_i;
  logic spi_flash_sd_3_o;
  logic spi_flash_sd_3_en_o;
  logic spi_flash_sd_3_i;
  modport ao_periph(
      input boot_select,
      input execute_from_flash,
      output exit_valid,
      output spi_flash_sck_o,
      output spi_flash_sck_en_o,
      output spi_flash_csb_0_o,
      output spi_flash_csb_0_en_o,
      output spi_flash_csb_1_o,
      output spi_flash_csb_1_en_o,
      output spi_flash_sd_0_o,
      output spi_flash_sd_0_en_o,
      input spi_flash_sd_0_i,
      output spi_flash_sd_1_o,
      output spi_flash_sd_1_en_o,
      input spi_flash_sd_1_i,
      output spi_flash_sd_2_o,
      output spi_flash_sd_2_en_o,
      input spi_flash_sd_2_i,
      output spi_flash_sd_3_o,
      output spi_flash_sd_3_en_o,
      input spi_flash_sd_3_i
  );
  modport pad_ring(
      output boot_select,
      output execute_from_flash,
      input exit_valid,
      input spi_flash_sck_o,
      input spi_flash_sck_en_o,
      input spi_flash_csb_0_o,
      input spi_flash_csb_0_en_o,
      input spi_flash_csb_1_o,
      input spi_flash_csb_1_en_o,
      input spi_flash_sd_0_o,
      input spi_flash_sd_0_en_o,
      output spi_flash_sd_0_i,
      input spi_flash_sd_1_o,
      input spi_flash_sd_1_en_o,
      output spi_flash_sd_1_i,
      input spi_flash_sd_2_o,
      input spi_flash_sd_2_en_o,
      output spi_flash_sd_2_i,
      input spi_flash_sd_3_o,
      input spi_flash_sd_3_en_o,
      output spi_flash_sd_3_i
  );
endinterface

interface if_bundle__ao_periph__core_v_mini_mcu ();
  logic rv_timer_0_intr;
  logic spi_flash_intr;
  logic rv_timer_1_intr;
  logic dma_done_intr;
  modport ao_periph(
      output rv_timer_0_intr,
      output spi_flash_intr,
      output rv_timer_1_intr,
      output dma_done_intr
  );
  modport core_v_mini_mcu(
      input rv_timer_0_intr,
      input spi_flash_intr,
      input rv_timer_1_intr,
      input dma_done_intr
  );
endinterface

interface if_bundle__pad_ring__pd_peripheral ();
  logic spi_host0_sd0_i;
  logic spi_host0_sd0_o;
  logic spi_host0_sd0_oe;
  logic spi_host0_sd1_i;
  logic spi_host0_sd1_o;
  logic spi_host0_sd1_oe;
  logic spi_host0_sd2_i;
  logic spi_host0_sd2_o;
  logic spi_host0_sd2_oe;
  logic spi_host0_sd3_i;
  logic spi_host0_sd3_o;
  logic spi_host0_sd3_oe;
  logic spi_host0_sck0_o;
  logic spi_host0_sck0_oe;
  logic spi_host0_csb0_o;
  logic spi_host0_csb0_oe;
  logic spi_host0_csb1_o;
  logic spi_host0_csb1_oe;
  logic io_pad_target_gpio_0_i;
  logic io_pad_target_gpio_0_o;
  logic io_pad_target_gpio_0_oe;
  logic io_pad_target_gpio_1_i;
  logic io_pad_target_gpio_1_o;
  logic io_pad_target_gpio_1_oe;
  logic io_pad_target_gpio_2_i;
  logic io_pad_target_gpio_2_o;
  logic io_pad_target_gpio_2_oe;
  logic io_pad_target_gpio_3_i;
  logic io_pad_target_gpio_3_o;
  logic io_pad_target_gpio_3_oe;
  logic io_pad_target_gpio_4_i;
  logic io_pad_target_gpio_4_o;
  logic io_pad_target_gpio_4_oe;
  logic io_pad_target_gpio_5_i;
  logic io_pad_target_gpio_5_o;
  logic io_pad_target_gpio_5_oe;
  logic io_pad_target_gpio_6_i;
  logic io_pad_target_gpio_6_o;
  logic io_pad_target_gpio_6_oe;
  logic io_pad_target_gpio_7_i;
  logic io_pad_target_gpio_7_o;
  logic io_pad_target_gpio_7_oe;
  logic io_pad_target_gpio_8_i;
  logic io_pad_target_gpio_8_o;
  logic io_pad_target_gpio_8_oe;
  logic io_pad_target_gpio_9_i;
  logic io_pad_target_gpio_9_o;
  logic io_pad_target_gpio_9_oe;
  logic io_pad_target_gpio_10_i;
  logic io_pad_target_gpio_10_o;
  logic io_pad_target_gpio_10_oe;
  logic io_pad_target_gpio_11_i;
  logic io_pad_target_gpio_11_o;
  logic io_pad_target_gpio_11_oe;
  logic io_pad_target_gpio_12_i;
  logic io_pad_target_gpio_12_o;
  logic io_pad_target_gpio_12_oe;
  logic io_pad_target_gpio_13_i;
  logic io_pad_target_gpio_13_o;
  logic io_pad_target_gpio_13_oe;
  logic io_pad_target_gpio_14_i;
  logic io_pad_target_gpio_14_o;
  logic io_pad_target_gpio_14_oe;
  logic io_pad_target_gpio_15_i;
  logic io_pad_target_gpio_15_o;
  logic io_pad_target_gpio_15_oe;
  logic io_pad_target_gpio_16_i;
  logic io_pad_target_gpio_16_o;
  logic io_pad_target_gpio_16_oe;
  logic io_pad_target_gpio_17_i;
  logic io_pad_target_gpio_17_o;
  logic io_pad_target_gpio_17_oe;
  logic uart0_rx0_i;
  logic uart0_tx0_o;
  logic uart0_tx0_oe;
  modport pd_peripheral(
      input spi_host0_sd0_i,
      output spi_host0_sd0_o,
      output spi_host0_sd0_oe,
      input spi_host0_sd1_i,
      output spi_host0_sd1_o,
      output spi_host0_sd1_oe,
      input spi_host0_sd2_i,
      output spi_host0_sd2_o,
      output spi_host0_sd2_oe,
      input spi_host0_sd3_i,
      output spi_host0_sd3_o,
      output spi_host0_sd3_oe,
      output spi_host0_sck0_o,
      output spi_host0_sck0_oe,
      output spi_host0_csb0_o,
      output spi_host0_csb0_oe,
      output spi_host0_csb1_o,
      output spi_host0_csb1_oe,
      input io_pad_target_gpio_0_i,
      output io_pad_target_gpio_0_o,
      output io_pad_target_gpio_0_oe,
      input io_pad_target_gpio_1_i,
      output io_pad_target_gpio_1_o,
      output io_pad_target_gpio_1_oe,
      input io_pad_target_gpio_2_i,
      output io_pad_target_gpio_2_o,
      output io_pad_target_gpio_2_oe,
      input io_pad_target_gpio_3_i,
      output io_pad_target_gpio_3_o,
      output io_pad_target_gpio_3_oe,
      input io_pad_target_gpio_4_i,
      output io_pad_target_gpio_4_o,
      output io_pad_target_gpio_4_oe,
      input io_pad_target_gpio_5_i,
      output io_pad_target_gpio_5_o,
      output io_pad_target_gpio_5_oe,
      input io_pad_target_gpio_6_i,
      output io_pad_target_gpio_6_o,
      output io_pad_target_gpio_6_oe,
      input io_pad_target_gpio_7_i,
      output io_pad_target_gpio_7_o,
      output io_pad_target_gpio_7_oe,
      input io_pad_target_gpio_8_i,
      output io_pad_target_gpio_8_o,
      output io_pad_target_gpio_8_oe,
      input io_pad_target_gpio_9_i,
      output io_pad_target_gpio_9_o,
      output io_pad_target_gpio_9_oe,
      input io_pad_target_gpio_10_i,
      output io_pad_target_gpio_10_o,
      output io_pad_target_gpio_10_oe,
      input io_pad_target_gpio_11_i,
      output io_pad_target_gpio_11_o,
      output io_pad_target_gpio_11_oe,
      input io_pad_target_gpio_12_i,
      output io_pad_target_gpio_12_o,
      output io_pad_target_gpio_12_oe,
      input io_pad_target_gpio_13_i,
      output io_pad_target_gpio_13_o,
      output io_pad_target_gpio_13_oe,
      input io_pad_target_gpio_14_i,
      output io_pad_target_gpio_14_o,
      output io_pad_target_gpio_14_oe,
      input io_pad_target_gpio_15_i,
      output io_pad_target_gpio_15_o,
      output io_pad_target_gpio_15_oe,
      input io_pad_target_gpio_16_i,
      output io_pad_target_gpio_16_o,
      output io_pad_target_gpio_16_oe,
      input io_pad_target_gpio_17_i,
      output io_pad_target_gpio_17_o,
      output io_pad_target_gpio_17_oe,
      input uart0_rx0_i,
      output uart0_tx0_o,
      output uart0_tx0_oe
  );
  modport pad_ring(
      output spi_host0_sd0_i,
      input spi_host0_sd0_o,
      input spi_host0_sd0_oe,
      output spi_host0_sd1_i,
      input spi_host0_sd1_o,
      input spi_host0_sd1_oe,
      output spi_host0_sd2_i,
      input spi_host0_sd2_o,
      input spi_host0_sd2_oe,
      output spi_host0_sd3_i,
      input spi_host0_sd3_o,
      input spi_host0_sd3_oe,
      input spi_host0_sck0_o,
      input spi_host0_sck0_oe,
      input spi_host0_csb0_o,
      input spi_host0_csb0_oe,
      input spi_host0_csb1_o,
      input spi_host0_csb1_oe,
      output io_pad_target_gpio_0_i,
      input io_pad_target_gpio_0_o,
      input io_pad_target_gpio_0_oe,
      output io_pad_target_gpio_1_i,
      input io_pad_target_gpio_1_o,
      input io_pad_target_gpio_1_oe,
      output io_pad_target_gpio_2_i,
      input io_pad_target_gpio_2_o,
      input io_pad_target_gpio_2_oe,
      output io_pad_target_gpio_3_i,
      input io_pad_target_gpio_3_o,
      input io_pad_target_gpio_3_oe,
      output io_pad_target_gpio_4_i,
      input io_pad_target_gpio_4_o,
      input io_pad_target_gpio_4_oe,
      output io_pad_target_gpio_5_i,
      input io_pad_target_gpio_5_o,
      input io_pad_target_gpio_5_oe,
      output io_pad_target_gpio_6_i,
      input io_pad_target_gpio_6_o,
      input io_pad_target_gpio_6_oe,
      output io_pad_target_gpio_7_i,
      input io_pad_target_gpio_7_o,
      input io_pad_target_gpio_7_oe,
      output io_pad_target_gpio_8_i,
      input io_pad_target_gpio_8_o,
      input io_pad_target_gpio_8_oe,
      output io_pad_target_gpio_9_i,
      input io_pad_target_gpio_9_o,
      input io_pad_target_gpio_9_oe,
      output io_pad_target_gpio_10_i,
      input io_pad_target_gpio_10_o,
      input io_pad_target_gpio_10_oe,
      output io_pad_target_gpio_11_i,
      input io_pad_target_gpio_11_o,
      input io_pad_target_gpio_11_oe,
      output io_pad_target_gpio_12_i,
      input io_pad_target_gpio_12_o,
      input io_pad_target_gpio_12_oe,
      output io_pad_target_gpio_13_i,
      input io_pad_target_gpio_13_o,
      input io_pad_target_gpio_13_oe,
      output io_pad_target_gpio_14_i,
      input io_pad_target_gpio_14_o,
      input io_pad_target_gpio_14_oe,
      output io_pad_target_gpio_15_i,
      input io_pad_target_gpio_15_o,
      input io_pad_target_gpio_15_oe,
      output io_pad_target_gpio_16_i,
      input io_pad_target_gpio_16_o,
      input io_pad_target_gpio_16_oe,
      output io_pad_target_gpio_17_i,
      input io_pad_target_gpio_17_o,
      input io_pad_target_gpio_17_oe,
      output uart0_rx0_i,
      input uart0_tx0_o,
      input uart0_tx0_oe
  );
endinterface

interface if_bundle__pd_peripheral__root ();
  logic spi_host1_sd0_i;
  logic spi_host1_sd0_o;
  logic spi_host1_sd0_oe;
  logic spi_host1_sd1_i;
  logic spi_host1_sd1_o;
  logic spi_host1_sd1_oe;
  logic spi_host1_sd2_i;
  logic spi_host1_sd2_o;
  logic spi_host1_sd2_oe;
  logic spi_host1_sd3_i;
  logic spi_host1_sd3_o;
  logic spi_host1_sd3_oe;
  logic spi_host1_sck0_o;
  logic spi_host1_sck0_oe;
  logic spi_host1_csb0_o;
  logic spi_host1_csb0_oe;
  logic spi_host1_csb1_o;
  logic spi_host1_csb1_oe;
  logic i2c0_sda0_i;
  logic i2c0_sda0_o;
  logic i2c0_sda0_oe;
  logic i2c0_scl0_i;
  logic i2c0_scl0_o;
  logic i2c0_scl0_oe;
  logic i2s0_sck0_i;
  logic i2s0_sck0_o;
  logic i2s0_sck0_oe;
  logic i2s0_ws0_i;
  logic i2s0_ws0_o;
  logic i2s0_ws0_oe;
  logic i2s0_sd0_i;
  logic i2s0_sd0_o;
  logic i2s0_sd0_oe;
  logic pdm2pcm0_pdm0_i;
  logic pdm2pcm0_pdm_clk0_o;
  logic io_pad_target_gpio_18_i;
  logic io_pad_target_gpio_18_o;
  logic io_pad_target_gpio_18_oe;
  logic io_pad_target_gpio_19_i;
  logic io_pad_target_gpio_19_o;
  logic io_pad_target_gpio_19_oe;
  logic io_pad_target_gpio_20_i;
  logic io_pad_target_gpio_20_o;
  logic io_pad_target_gpio_20_oe;
  logic io_pad_target_gpio_21_i;
  logic io_pad_target_gpio_21_o;
  logic io_pad_target_gpio_21_oe;
  logic io_pad_target_gpio_22_i;
  logic io_pad_target_gpio_22_o;
  logic io_pad_target_gpio_22_oe;
  logic io_pad_target_gpio_23_i;
  logic io_pad_target_gpio_23_o;
  logic io_pad_target_gpio_23_oe;
  logic io_pad_target_gpio_24_i;
  logic io_pad_target_gpio_24_o;
  logic io_pad_target_gpio_24_oe;
  logic io_pad_target_gpio_25_i;
  logic io_pad_target_gpio_25_o;
  logic io_pad_target_gpio_25_oe;
  logic io_pad_target_gpio_26_i;
  logic io_pad_target_gpio_26_o;
  logic io_pad_target_gpio_26_oe;
  logic io_pad_target_gpio_27_i;
  logic io_pad_target_gpio_27_o;
  logic io_pad_target_gpio_27_oe;
  logic io_pad_target_gpio_28_i;
  logic io_pad_target_gpio_28_o;
  logic io_pad_target_gpio_28_oe;
  logic io_pad_target_gpio_29_i;
  logic io_pad_target_gpio_29_o;
  logic io_pad_target_gpio_29_oe;
  logic io_pad_target_gpio_30_i;
  logic io_pad_target_gpio_30_o;
  logic io_pad_target_gpio_30_oe;
  logic io_pad_target_gpio_31_i;
  logic io_pad_target_gpio_31_o;
  logic io_pad_target_gpio_31_oe;
  logic ext_intr_0;
  logic ext_intr_1;
  modport pd_peripheral(
      input spi_host1_sd0_i,
      output spi_host1_sd0_o,
      output spi_host1_sd0_oe,
      input spi_host1_sd1_i,
      output spi_host1_sd1_o,
      output spi_host1_sd1_oe,
      input spi_host1_sd2_i,
      output spi_host1_sd2_o,
      output spi_host1_sd2_oe,
      input spi_host1_sd3_i,
      output spi_host1_sd3_o,
      output spi_host1_sd3_oe,
      output spi_host1_sck0_o,
      output spi_host1_sck0_oe,
      output spi_host1_csb0_o,
      output spi_host1_csb0_oe,
      output spi_host1_csb1_o,
      output spi_host1_csb1_oe,
      input i2c0_sda0_i,
      output i2c0_sda0_o,
      output i2c0_sda0_oe,
      input i2c0_scl0_i,
      output i2c0_scl0_o,
      output i2c0_scl0_oe,
      input i2s0_sck0_i,
      output i2s0_sck0_o,
      output i2s0_sck0_oe,
      input i2s0_ws0_i,
      output i2s0_ws0_o,
      output i2s0_ws0_oe,
      input i2s0_sd0_i,
      output i2s0_sd0_o,
      output i2s0_sd0_oe,
      input pdm2pcm0_pdm0_i,
      output pdm2pcm0_pdm_clk0_o,
      input io_pad_target_gpio_18_i,
      output io_pad_target_gpio_18_o,
      output io_pad_target_gpio_18_oe,
      input io_pad_target_gpio_19_i,
      output io_pad_target_gpio_19_o,
      output io_pad_target_gpio_19_oe,
      input io_pad_target_gpio_20_i,
      output io_pad_target_gpio_20_o,
      output io_pad_target_gpio_20_oe,
      input io_pad_target_gpio_21_i,
      output io_pad_target_gpio_21_o,
      output io_pad_target_gpio_21_oe,
      input io_pad_target_gpio_22_i,
      output io_pad_target_gpio_22_o,
      output io_pad_target_gpio_22_oe,
      input io_pad_target_gpio_23_i,
      output io_pad_target_gpio_23_o,
      output io_pad_target_gpio_23_oe,
      input io_pad_target_gpio_24_i,
      output io_pad_target_gpio_24_o,
      output io_pad_target_gpio_24_oe,
      input io_pad_target_gpio_25_i,
      output io_pad_target_gpio_25_o,
      output io_pad_target_gpio_25_oe,
      input io_pad_target_gpio_26_i,
      output io_pad_target_gpio_26_o,
      output io_pad_target_gpio_26_oe,
      input io_pad_target_gpio_27_i,
      output io_pad_target_gpio_27_o,
      output io_pad_target_gpio_27_oe,
      input io_pad_target_gpio_28_i,
      output io_pad_target_gpio_28_o,
      output io_pad_target_gpio_28_oe,
      input io_pad_target_gpio_29_i,
      output io_pad_target_gpio_29_o,
      output io_pad_target_gpio_29_oe,
      input io_pad_target_gpio_30_i,
      output io_pad_target_gpio_30_o,
      output io_pad_target_gpio_30_oe,
      input io_pad_target_gpio_31_i,
      output io_pad_target_gpio_31_o,
      output io_pad_target_gpio_31_oe,
      input ext_intr_0,
      input ext_intr_1
  );
  modport root(
      output spi_host1_sd0_i,
      input spi_host1_sd0_o,
      input spi_host1_sd0_oe,
      output spi_host1_sd1_i,
      input spi_host1_sd1_o,
      input spi_host1_sd1_oe,
      output spi_host1_sd2_i,
      input spi_host1_sd2_o,
      input spi_host1_sd2_oe,
      output spi_host1_sd3_i,
      input spi_host1_sd3_o,
      input spi_host1_sd3_oe,
      input spi_host1_sck0_o,
      input spi_host1_sck0_oe,
      input spi_host1_csb0_o,
      input spi_host1_csb0_oe,
      input spi_host1_csb1_o,
      input spi_host1_csb1_oe,
      output i2c0_sda0_i,
      input i2c0_sda0_o,
      input i2c0_sda0_oe,
      output i2c0_scl0_i,
      input i2c0_scl0_o,
      input i2c0_scl0_oe,
      output i2s0_sck0_i,
      input i2s0_sck0_o,
      input i2s0_sck0_oe,
      output i2s0_ws0_i,
      input i2s0_ws0_o,
      input i2s0_ws0_oe,
      output i2s0_sd0_i,
      input i2s0_sd0_o,
      input i2s0_sd0_oe,
      output pdm2pcm0_pdm0_i,
      input pdm2pcm0_pdm_clk0_o,
      output io_pad_target_gpio_18_i,
      input io_pad_target_gpio_18_o,
      input io_pad_target_gpio_18_oe,
      output io_pad_target_gpio_19_i,
      input io_pad_target_gpio_19_o,
      input io_pad_target_gpio_19_oe,
      output io_pad_target_gpio_20_i,
      input io_pad_target_gpio_20_o,
      input io_pad_target_gpio_20_oe,
      output io_pad_target_gpio_21_i,
      input io_pad_target_gpio_21_o,
      input io_pad_target_gpio_21_oe,
      output io_pad_target_gpio_22_i,
      input io_pad_target_gpio_22_o,
      input io_pad_target_gpio_22_oe,
      output io_pad_target_gpio_23_i,
      input io_pad_target_gpio_23_o,
      input io_pad_target_gpio_23_oe,
      output io_pad_target_gpio_24_i,
      input io_pad_target_gpio_24_o,
      input io_pad_target_gpio_24_oe,
      output io_pad_target_gpio_25_i,
      input io_pad_target_gpio_25_o,
      input io_pad_target_gpio_25_oe,
      output io_pad_target_gpio_26_i,
      input io_pad_target_gpio_26_o,
      input io_pad_target_gpio_26_oe,
      output io_pad_target_gpio_27_i,
      input io_pad_target_gpio_27_o,
      input io_pad_target_gpio_27_oe,
      output io_pad_target_gpio_28_i,
      input io_pad_target_gpio_28_o,
      input io_pad_target_gpio_28_oe,
      output io_pad_target_gpio_29_i,
      input io_pad_target_gpio_29_o,
      input io_pad_target_gpio_29_oe,
      output io_pad_target_gpio_30_i,
      input io_pad_target_gpio_30_o,
      input io_pad_target_gpio_30_oe,
      output io_pad_target_gpio_31_i,
      input io_pad_target_gpio_31_o,
      input io_pad_target_gpio_31_oe,
      output ext_intr_0,
      output ext_intr_1
  );
endinterface

interface if_bundle__core_v_mini_mcu__pd_peripheral ();
  logic rv_plic_0_irq;
  logic rv_plic_0_msip;
  logic rv_timer_2_3_timer_expired_0_0_intr_o;
  logic rv_timer_2_3_timer_expired_1_0_intr_o;
  logic spi_host_0_spi_event_intr_o;
  logic gpio_0_intr_o;
  logic gpio_1_intr_o;
  logic gpio_2_intr_o;
  logic gpio_3_intr_o;
  logic gpio_4_intr_o;
  logic gpio_5_intr_o;
  logic gpio_6_intr_o;
  logic gpio_7_intr_o;
  modport pd_peripheral(
      output rv_plic_0_irq,
      output rv_plic_0_msip,
      output rv_timer_2_3_timer_expired_0_0_intr_o,
      output rv_timer_2_3_timer_expired_1_0_intr_o,
      output spi_host_0_spi_event_intr_o,
      output gpio_0_intr_o,
      output gpio_1_intr_o,
      output gpio_2_intr_o,
      output gpio_3_intr_o,
      output gpio_4_intr_o,
      output gpio_5_intr_o,
      output gpio_6_intr_o,
      output gpio_7_intr_o
  );
  modport core_v_mini_mcu(
      input rv_plic_0_irq,
      input rv_plic_0_msip,
      input rv_timer_2_3_timer_expired_0_0_intr_o,
      input rv_timer_2_3_timer_expired_1_0_intr_o,
      input spi_host_0_spi_event_intr_o,
      input gpio_0_intr_o,
      input gpio_1_intr_o,
      input gpio_2_intr_o,
      input gpio_3_intr_o,
      input gpio_4_intr_o,
      input gpio_5_intr_o,
      input gpio_6_intr_o,
      input gpio_7_intr_o
  );
endinterface

interface if_bundle__ao_periph__root ();
  logic dma_ext_rx;
  logic dma_ext_tx;
  modport root(output dma_ext_rx, output dma_ext_tx);
  modport ao_periph(input dma_ext_rx, input dma_ext_tx);
endinterface

interface if_bundle__ao_periph__pd_peripheral ();
  logic dma_window_intr;
  logic spi_host_0_rx_valid;
  logic spi_host_0_tx_valid;
  logic i2s_0_rx_valid;
  modport ao_periph(
      output dma_window_intr,
      input spi_host_0_rx_valid,
      input spi_host_0_tx_valid,
      input i2s_0_rx_valid
  );
  modport pd_peripheral(
      input dma_window_intr,
      output spi_host_0_rx_valid,
      output spi_host_0_tx_valid,
      output i2s_0_rx_valid
  );
endinterface


/* verilator lint_on DECLFILENAME */
