// Copyright EPFL contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

module myinverter (
    input  logic a,
    output logic z
);

endmodule : myinverter

