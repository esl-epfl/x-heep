// Copyright 2018 Robert Balas <balasr@student.ethz.ch>
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Contributor: Robert Balas <balasr@student.ethz.ch>

module core_v_mini_mcu #(
    parameter PULP_XPULP = 0,
    parameter FPU        = 0,
    parameter PULP_ZFINX = 0
) (
    input logic clk_i,
    input logic rst_ni,

    input  logic        jtag_tck_i,
    input  logic        jtag_tms_i,
    input  logic        jtag_trst_ni,
    input  logic        jtag_tdi_i,
    output logic        jtag_tdo_o,

    input  logic        fetch_enable_i,
    output logic [31:0] exit_value_o,
    output logic        exit_valid_o
);

  `include "tb_util.svh"

  import core_v_mini_mcu_pkg::*;
  import obi_pkg::*;
  import cv32e40p_apu_core_pkg::*;

  localparam NUM_BYTES      = 2**16; //must be 2**16, it is not a parameter!!!
  localparam DM_HALTADDRESS = core_v_mini_mcu_pkg::DEBUG_START_ADDRESS + 32'h00000800; //debug rom code (section .text in linker) starts at 0x800

  localparam JTAG_IDCODE      = 32'h10001c05;
  localparam BOOT_ADDR        = 'h180;
  localparam NUM_MHPMCOUNTERS = 1;


  // signals connecting core to memory

  obi_req_t     core_instr_req;
  obi_resp_t    core_instr_resp;
  obi_req_t     core_data_req;
  obi_resp_t    core_data_resp;
  obi_req_t     debug_master_req;
  obi_resp_t    debug_master_resp;

  obi_req_t     ram0_slave_req;
  obi_resp_t    ram0_slave_resp;
  obi_req_t     ram1_slave_req;
  obi_resp_t    ram1_slave_resp;
  obi_req_t     debug_slave_req;
  obi_resp_t    debug_slave_resp;
  obi_req_t     peripheral_slave_req;
  obi_resp_t    peripheral_slave_resp;

  // signals to debug unit
  logic                               debug_core_req;

  // irq signals
  logic                               irq_ack;
  logic [                  4:0]       irq_id_out;
  logic                               irq_software;
  logic                               irq_timer;
  logic                               irq_external;
  logic [                 15:0]       irq_fast;


  cpu_subsystem #(
    .BOOT_ADDR        (BOOT_ADDR),
    .PULP_XPULP       (PULP_XPULP),
    .FPU              (FPU),
    .PULP_ZFINX       (PULP_ZFINX),
    .NUM_MHPMCOUNTERS (NUM_MHPMCOUNTERS),
    .DM_HALTADDRESS   (DM_HALTADDRESS)
  ) cpu_subsystem_i (
      // Clock and Reset
      .clk_i,
      .rst_ni,
      .core_instr_req_o(core_instr_req),
      .core_instr_resp_i(core_instr_resp),
      .core_data_req_o(core_data_req),
      .core_data_resp_i(core_data_resp),
      .irq_i({irq_fast, 4'b0, irq_external, 3'b0, irq_timer, 3'b0, irq_software, 3'b0}),
      .irq_ack_o(irq_ack),
      .irq_id_o(irq_id_out),
      .debug_req_i(debug_core_req),
      .fetch_enable_i(fetch_enable_i)
  );


  debug_subsystem #(
      .JTAG_IDCODE(JTAG_IDCODE)
  ) debug_subsystem_i (
    .clk_i               ( clk_i            ),
    .rst_ni              ( rst_ni           ),

    .jtag_tck_i          ( jtag_tck_i       ),
    .jtag_tms_i          ( jtag_tms_i       ),
    .jtag_trst_ni        ( jtag_trst_ni     ),
    .jtag_tdi_i          ( jtag_tdi_i       ),
    .jtag_tdo_o          ( jtag_tdo_o       ),

    .debug_core_req_o    ( debug_core_req   ),

    .debug_slave_req_i   ( debug_slave_req   ),
    .debug_slave_resp_o  ( debug_slave_resp  ),
    .debug_master_req_o  ( debug_master_req  ),
    .debug_master_resp_i ( debug_master_resp )

  );

  system_bus #(
      .NUM_BYTES(NUM_BYTES)
  ) system_bus_i (
    .clk_i (clk_i),
    .rst_ni(rst_ni),

    .core_instr_req_i        ( core_instr_req        ),
    .core_instr_resp_o       ( core_instr_resp       ),
    .core_data_req_i         ( core_data_req         ),
    .core_data_resp_o        ( core_data_resp        ),
    .debug_master_req_i      ( debug_master_req      ),
    .debug_master_resp_o     ( debug_master_resp     ),

    .ram0_req_o              ( ram0_slave_req        ),
    .ram0_resp_i             ( ram0_slave_resp       ),
    .ram1_req_o              ( ram1_slave_req        ),
    .ram1_resp_i             ( ram1_slave_resp       ),
    .debug_slave_req_o       ( debug_slave_req       ),
    .debug_slave_resp_i      ( debug_slave_resp      ),
    .peripheral_slave_req_o  ( peripheral_slave_req  ),
    .peripheral_slave_resp_i ( peripheral_slave_resp )

  );

  memory_subsystem #(
      .NUM_BYTES(NUM_BYTES)
  ) memory_subsystem_i (
    .clk_i,
    .rst_ni,
    .ram0_req_i(ram0_slave_req),
    .ram0_resp_o(ram0_slave_resp),
    .ram1_req_i(ram1_slave_req),
    .ram1_resp_o(ram1_slave_resp)
  );

  peripheral_subsystem peripheral_subsystem_i
  (
    .clk_i,
    .rst_ni,

    .slave_req_i(peripheral_slave_req),
    .slave_resp_o(peripheral_slave_resp),

    .exit_valid_o  (exit_valid_o),
    .exit_value_o  (exit_value_o),

    .uart_rx_i('0),
    .uart_tx_o(),
    .uart_tx_en_o(),
    .uart_intr_tx_watermark_o() ,
    .uart_intr_rx_watermark_o() ,
    .uart_intr_tx_empty_o()  ,
    .uart_intr_rx_overflow_o()  ,
    .uart_intr_rx_frame_err_o() ,
    .uart_intr_rx_break_err_o() ,
    .uart_intr_rx_timeout_o()   ,
    .uart_intr_rx_parity_err_o()
  );

  assign irq_software = '0;
  assign irq_timer    = '0;
  assign irq_external = '0;
  assign irq_fast     = '0;


endmodule  // cv32e40p_tb_subsystem
