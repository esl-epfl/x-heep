/*
 * Copyright 2025 EPFL
 * Solderpad Hardware License, Version 2.1, see LICENSE.md for details.
 * SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 *
 * Author: Tommaso Terzano <tommaso.terzano@epfl.ch>
 *                         <tommaso.terzano@gmail.com>
 *
 * Info: Header file for the DMA subsystem.
 */



`define ADDR_MODE_EN
`define ZERO_PADDING_EN
`define SUBADDR_MODE_EN
`define HW_FIFO_MODE_EN
